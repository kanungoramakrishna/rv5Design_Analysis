import rv32i_types::*;
import alumux::*;
import cmpmux::*;

module ex_forward_unit 
(
	// TODO I/O
);

// TODO implement

endmodule 