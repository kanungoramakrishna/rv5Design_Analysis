import rv32i_types::*;

module mem_forward_unit
(
	// TODO I/O
);

// TODO implement

endmodule
