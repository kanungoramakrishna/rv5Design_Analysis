module memory_access
(

);