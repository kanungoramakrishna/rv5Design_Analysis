import rv32i_types::*;

module hazard_unit
(
	// TODO I/O
);

// TODO implement

endmodule