import rv32i_types::*;

module branch_predictor
(
	// TODO
);

// TODO

endmodule