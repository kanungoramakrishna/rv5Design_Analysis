module execute
(

);