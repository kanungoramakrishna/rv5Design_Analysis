module write_back
(

);