module instruction_fetch
(

);